module data_memory #(
    parameter W=`WORD_WIDTH
) (
    input clk,rst,
    
);
    
endmodule